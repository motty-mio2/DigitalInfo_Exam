module PENC4(A, Y, VALID); // A：4 bit 入力，Y：2 bit エンコード出力，VALID：有効信号（= 1：Y 出力有効）
endmodule